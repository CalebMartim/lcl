module exp(
	
);
endmodule
